`timescale 1ns / 1ps


module inst_mem(Address, Instruction); 

    input [7:0] Address; 

    output [15:0] Instruction;
    
    reg [15:0] mem[0:32];

	initial
	begin
		mem[8'h00] = 16'b0000000100101111;
		mem[8'h02] = 16'b0000000100101110;
		mem[8'h04] = 16'b0000001101001100;
		mem[8'h06] = 16'b0000001100101101;
		
		mem[8'h08] = 16'b0000010101100001;
		mem[8'h0a] = 16'b0000000101010010;
		mem[8'h0c] = 16'b0000000000001110;
		mem[8'h0e] = 16'b0000010000111010;
		
		mem[8'h10] = 16'b0000010000101011;
		mem[8'h12] = 16'b0000011000111001;
		mem[8'h14] = 16'b0000011000101000;
		mem[8'h16] = 16'b0110011100001100;
		
		mem[8'h18] = 16'b0000101100011111;
		mem[8'h1a] = 16'b0100011100001101;
		mem[8'h1c] = 16'b0000101100101111;
		mem[8'h1e] = 16'b0101010000001010;
		
		mem[8'h20] = 16'b0000000100011111;
		mem[8'h22] = 16'b0000000100011111;
		mem[8'h24] = 16'b1000100000001001;
		mem[8'h26] = 16'b0000100010001111;
		
		mem[8'h28] = 16'b1011100000101001;
		mem[8'h2a] = 16'b1000101000101001;
		mem[8'h2c] = 16'b0000110011001111;
		mem[8'h2e] = 16'b0000110111011110;
		
		mem[8'h30] = 16'b0000110011011111;
		mem[8'h32] = 16'b1110111111111111;
		mem[8'h34] = 16'b0000000000000000;
		mem[8'h36] = 16'b0000000000000000;
		
		mem[8'h38] = 16'b0000000000000000;
		mem[8'h3a] = 16'b0000000000000000;
		mem[8'h3c] = 16'b0000000000000000;
		mem[8'h3e] = 16'b0000000000000000;
		
	end

	assign Instruction = mem[Address];	
	

endmodule