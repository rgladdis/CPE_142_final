module shift_left1(a, y);

input a;
output y;

assign y = a << 1;

endmodule